`include "bsg_defines.v"

`include "bsg_clk_gen.vh"

module bsg_dmc_clk_rst_gen
  import bsg_tag_pkg::bsg_tag_s;
  import bsg_dmc_pkg::*;
 #(parameter num_adgs_p         = 2
  ,parameter `BSG_INV_PARAM(dq_group_p        ))
  (
  input bsg_dmc_dly_tag_lines_s    dly_tag_lines_i
  ,input bsg_dmc_osc_tag_lines_s     osc_tag_lines_i    
  // asynchronous reset for dram controller
  ,output                            async_reset_o
  // clock input and delayed clock output (for dqs), generating 90-degree phase
  // shift
  ,input            [dq_group_p-1:0] dqs_clk_i
  ,output           [dq_group_p-1:0] dqs_clk_o
  // 2x clock input from clock generator and 1x clock output
  ,input                             ext_dfi_clk_2x_i
  ,output                            dfi_clk_2x_o
  ,output                            dfi_clk_1x_o
  ,output							 clock_monitor_clk_o);

  localparam debug_level_lp = 0;

  genvar i;

  bsg_tag_client_unsync #(.width_p(1)) btc_async_reset
    (.bsg_tag_i      ( dly_tag_lines_i.async_reset_tag )
    ,.data_async_r_o ( async_reset_o     ));

  // Clock Generator (CG) Instance
  for(i=0;i<dq_group_p;i++) begin: dly_lines
    bsg_dly_line #(.num_adgs_p(num_adgs_p)) dly_line_inst
      (.bsg_tag_i         ( dly_tag_lines_i.bsg_dly_tag[i]         )
      ,.bsg_tag_trigger_i ( dly_tag_lines_i.bsg_dly_trigger_tag[i] )
      ,.async_reset_i     ( async_reset_o            )
      ,.clk_i             ( dqs_clk_i[i]             )
      ,.clk_o             ( dqs_clk_o[i]             ));
  end

  `declare_bsg_clk_gen_ds_tag_payload_s(2)

  bsg_clk_gen_ds_tag_payload_s ds_tag_payload_r;

  bsg_clk_gen_ds_tag_payload_s clk_monitor_ds_tag_payload_r;

  wire  ds_tag_payload_new_r;

  // fixme: maybe wire up a default and deal with reset issue?
  // downsampler bsg_tag interface
  bsg_tag_client #
    (.width_p   ( $bits(bsg_clk_gen_ds_tag_payload_s) )
    ,.harden_p  ( 1                                   ))
  btc_ds
    (.bsg_tag_i     ( dly_tag_lines_i.bsg_ds_tag         )

    ,.recv_clk_i    ( dfi_clk_2x_o             )
    ,.recv_new_r_o  ( ds_tag_payload_new_r )   // we don't require notification
    ,.recv_data_r_o ( ds_tag_payload_r     ));

  bsg_tag_client #
    (.width_p   ( $bits(bsg_clk_gen_ds_tag_payload_s) )
    ,.harden_p  ( 1                                   ))
  btc_clk_monitor_ds
    (.bsg_tag_i     (osc_tag_lines_i.bsg_clk_monitor_ds_tag)

    ,.recv_clk_i    ( dfi_clk_2x_o             )
    ,.recv_new_r_o  (  )   // we don't require notification
    ,.recv_data_r_o ( clk_monitor_ds_tag_payload_r     ));


  // synopsys translate_off
  if (debug_level_lp > 1)
  always_ff @(negedge dfi_clk_2x_o) begin
    if (ds_tag_payload_new_r)
      $display("## bsg_clk_gen downsampler received configuration state: %b",ds_tag_payload_r);
  end
  // synopsys translate_on

  // clock downsampler
  //
  // we allow the clock downsample reset to be accessed via bsg_tag; this way
  // we can turn it off by holding reset high to save power.
  //
  bsg_counter_clock_downsample #
    (.width_p  ( 2 )
    ,.harden_p ( 1 ))
  clk_gen_ds_inst
    (.clk_i   ( dfi_clk_2x_o           )
    ,.reset_i ( ds_tag_payload_r.reset )
    ,.val_i   ( 2'd0                   ) // Always 2X->1X
    ,.clk_r_o ( dfi_clk_1x_o           ));

  bsg_counter_clock_downsample #
    (.width_p  ( 2 )
    ,.harden_p ( 1 ))
  clk_monitor_clk_gen
    (.clk_i   ( dfi_clk_2x_o               )
    ,.reset_i ( clk_monitor_ds_tag_payload_r.reset )
    ,.val_i   ( clk_monitor_ds_tag_payload_r.val )
    //,.val_i   ( 2'b1 )	
    ,.clk_r_o (clock_monitor_clk_o	   ));

  logic async_reset_lo;

  bsg_tag_client_unsync #( .width_p(1) )
    osc_async_reset
      (.bsg_tag_i(osc_tag_lines_i.async_reset)
      ,.data_async_r_o(async_reset_lo)
      );

  bsg_clk_gen #(.downsample_width_p(2)
               ,.num_adgs_p(num_adgs_p)
               ,.version_p(2)
  			 ,.nonsynth_sim_osc_granularity_p(50)
               )
  clk_gen_inst
      (.async_osc_reset_i     (async_reset_lo)
      ,.bsg_osc_tag_i         (osc_tag_lines_i.osc)
      ,.bsg_osc_trigger_tag_i (osc_tag_lines_i.osc_trigger)
      ,.bsg_ds_tag_i          (osc_tag_lines_i.ds)
      ,.ext_clk_i             (ext_dfi_clk_2x_i)
      ,.select_i              (osc_tag_lines_i.sel)
      ,.clk_o                 (dfi_clk_2x_o)
      );

endmodule

`BSG_ABSTRACT_MODULE(bsg_dmc_clk_rst_gen)
